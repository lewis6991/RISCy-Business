//----------------------------------------
// File: ex_control_tb.sv
// Description: Execute controller testbench
// Primary Author: Jack Barnes
// Other Contributors:
// Notes: Full test coverage
//----------------------------------------
module ex_control_tb;

timeunit 10ns; timeprecision 100ps;
const int clk = 100;

ex_control ex_control0 (
);

//Initial conditions
initial
begin
end

//Testing procedure
initial
begin
end

endmodule
