//----------------------------------------
// File: alu_tb.sv
// Description: PC testbench
// Primary Author: Jack Barnes
// Other Contributors:
// Notes: Full test coverage of ALU instructions
//        Select sample for each instruction
//----------------------------------------
module alu_tb;

timeunit 10ns; timeprecision 100ps;
const int clk = 100;

alu alu0 (
);

//Initial conditions
initial
begin
end

//Testing procedure
initial
begin
end

endmodule
