//----------------------------------------
// File: decoder_t.sv
// Description: Decoder testbench
// Primary Author: Jack
// Other Contributors:
// Notes: Full test coverage
//----------------------------------------
module decoder_t;

const int clk = 100;

decoder decoder0 (
);

//Initial conditions
initial
begin
end

//Testing procedure
initial
begin
end

endmodule
