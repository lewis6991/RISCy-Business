//------------------------------------------------------------------------------
// File              : ex_mult.sv
// Description       : MULT module for execute stage
// Primary Author    : Ethan Bishop
// Other Contributors:
// Notes             :
//------------------------------------------------------------------------------
module ex_mult (
    input        [31:0] A     ,
                        B     ,
    input               SelB  , // Enable B input, else multiply by 1
    input        [5:0]  OpCode,
                        Func  ,
    output logic        C     ,
                        Z     ,
                        O     ,
                        N     ,
    output logic [63:0] Out   ,
    output logic [31:0] mB
);

    always_comb
    begin
        mB = SelB ? B : 32'd1;

        case (Func)
            `CLZ:
                casez (A)
                    32'b1???????????????????????????????: Out = 0 ;
                    32'b01??????????????????????????????: Out = 1 ;
                    32'b001?????????????????????????????: Out = 2 ;
                    32'b0001????????????????????????????: Out = 3 ;
                    32'b00001???????????????????????????: Out = 4 ;
                    32'b000001??????????????????????????: Out = 5 ;
                    32'b0000001?????????????????????????: Out = 6 ;
                    32'b00000001????????????????????????: Out = 7 ;
                    32'b000000001???????????????????????: Out = 8 ;
                    32'b0000000001??????????????????????: Out = 9 ;
                    32'b00000000001?????????????????????: Out = 10;
                    32'b000000000001????????????????????: Out = 11;
                    32'b0000000000001???????????????????: Out = 12;
                    32'b00000000000001??????????????????: Out = 13;
                    32'b000000000000001?????????????????: Out = 14;
                    32'b0000000000000001????????????????: Out = 15;
                    32'b00000000000000001???????????????: Out = 16;
                    32'b000000000000000001??????????????: Out = 17;
                    32'b0000000000000000001?????????????: Out = 18;
                    32'b00000000000000000001????????????: Out = 19;
                    32'b000000000000000000001???????????: Out = 20;
                    32'b0000000000000000000001??????????: Out = 21;
                    32'b00000000000000000000001?????????: Out = 22;
                    32'b000000000000000000000001????????: Out = 23;
                    32'b0000000000000000000000001???????: Out = 24;
                    32'b00000000000000000000000001??????: Out = 25;
                    32'b000000000000000000000000001?????: Out = 26;
                    32'b0000000000000000000000000001????: Out = 27;
                    32'b00000000000000000000000000001???: Out = 28;
                    32'b000000000000000000000000000001??: Out = 29;
                    32'b0000000000000000000000000000001?: Out = 30;
                    32'b00000000000000000000000000000001: Out = 31;
                    32'b00000000000000000000000000000000: Out = 32;
                endcase
            `CLO:
                casez (A)
                    32'b0???????????????????????????????: Out = 0 ;
                    32'b10??????????????????????????????: Out = 1 ;
                    32'b110?????????????????????????????: Out = 2 ;
                    32'b1110????????????????????????????: Out = 3 ;
                    32'b11110???????????????????????????: Out = 4 ;
                    32'b111110??????????????????????????: Out = 5 ;
                    32'b1111110?????????????????????????: Out = 6 ;
                    32'b11111110????????????????????????: Out = 7 ;
                    32'b111111110???????????????????????: Out = 8 ;
                    32'b1111111110??????????????????????: Out = 9 ;
                    32'b11111111110?????????????????????: Out = 10;
                    32'b111111111110????????????????????: Out = 11;
                    32'b1111111111110???????????????????: Out = 12;
                    32'b11111111111110??????????????????: Out = 13;
                    32'b111111111111110?????????????????: Out = 14;
                    32'b1111111111111110????????????????: Out = 15;
                    32'b11111111111111110???????????????: Out = 16;
                    32'b111111111111111110??????????????: Out = 17;
                    32'b1111111111111111110?????????????: Out = 18;
                    32'b11111111111111111110????????????: Out = 19;
                    32'b111111111111111111110???????????: Out = 20;
                    32'b1111111111111111111110??????????: Out = 21;
                    32'b11111111111111111111110?????????: Out = 22;
                    32'b111111111111111111111110????????: Out = 23;
                    32'b1111111111111111111111110???????: Out = 24;
                    32'b11111111111111111111111110??????: Out = 25;
                    32'b111111111111111111111111110?????: Out = 26;
                    32'b1111111111111111111111111110????: Out = 27;
                    32'b11111111111111111111111111110???: Out = 28;
                    32'b111111111111111111111111111110??: Out = 29;
                    32'b1111111111111111111111111111110?: Out = 31;
                    32'b11111111111111111111111111111110: Out = 31;
                    32'b11111111111111111111111111111111: Out = 32;
                endcase
                default: Out = A;
        endcase

        C = Out[32]       ;
        Z = Out[31:0] == 0;
        O = Out[32]       ;
        N = Out[31]       ;

    end

endmodule
