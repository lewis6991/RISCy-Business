//------------------------------------------------------------------------------
// File              : Control.sv
// Description       : Control module.
// Author            :
// Other Contributers:
// Notes             :
//------------------------------------------------------------------------------

module control(
    input Clock ,
    input nReset,
);

endmodule
