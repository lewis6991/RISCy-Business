//----------------------------------------
// File: decoder_tb.sv
// Description: Decoder testbench
// Primary Author: Jack Barnes
// Other Contributors:
// Notes: Full test coverage
//----------------------------------------
module decoder_tb;

timeunit 10ns; timeprecision 100ps;
const int clk = 100;

decoder decoder0 (
);

//Initial conditions
initial
begin
end

//Testing procedure
initial
begin
end

endmodule
