//----------------------------------------
// File: IF_tb.sv
// Description: Instruction Fetch testbench
// Primary Author: Jack Barnes
// Other Contributors:
// Notes: Full test coverage
//----------------------------------------
module IF_tb;

timeunit 10ns; timeprecision 100ps;
const int clk = 100;

IF IF0 (
);

//Initial conditions
initial
begin
end

//Testing procedure
initial
begin
end

endmodule
