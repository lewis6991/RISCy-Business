/------------------------------------------------------------------------------
// File              : BP.sv
// Description       : Branch prediction unit
// Primary Author    : -
// Other Contributors: 
// Notes             : Placeholder
//------------------------------------------------------------------------------

module BP(
);

endmodule
