//------------------------------------------------------------------------------
// File              : processor.sv
// Description       : Top-level module for MIPS32 processor.
// Primary Author    :
// Other Contributers: Lewis Russell
// Notes             :
//------------------------------------------------------------------------------

module processor(
    input logic Clock,
    input logic nReset
);

endmodule
