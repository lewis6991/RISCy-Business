//------------------------------------------------------------------------------
// File              : mem_func.sv
// Description       : Memory Functions Codes (Extracted from Opcode)
// Primary Author    : Dhanushan Raveendran
// Other Contributors: 
// Notes             :  
//------------------------------------------------------------------------------

`define BS 3'b000
`define BU 3'b100
`define HS 3'b001
`define HU 3'b101
`define WD 3'b011
`define WL 3'b010
`define WR 3'b110
