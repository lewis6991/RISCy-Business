//----------------------------------------
// File: mul_definition.sv
// Description: MUL instruction codes
// Primary Author: Dhanushan
// Other Contributors: 
// Notes: 
//----------------------------------------

`define		CLO		6'b100001
`define		CLZ		6'b100000

`define		MADD	6'b000000
`define		MADDU	6'b000001
`define		MSUB	6'b000100
`define		MSUBU	6'b000101
`define		MUL		6'b000010	