//----------------------------------------
// File: alu_t.sv
// Description: PC testbench
// Primary Author: Jack
// Other Contributors:
// Notes: Full test coverage of ALU instructions
//        Select sample for each instruction
//----------------------------------------
module alu_t;

const int clk = 100;

alu alu0 (
);

//Initial conditions
initial
begin
end

//Testing procedure
initial
begin
end

endmodule
