//----------------------------------------
// File: BP_tb.sv
// Description: Branch prediction testbench
// Primary Author: Jack Barnes
// Other Contributors:
// Notes: Full test coverage
//----------------------------------------
module BP_tb;

timeunit 10ns; timeprecision 100ps;
const int clk = 100;

BP BP0 (
);

//Initial conditions
initial
begin
end

//Testing procedure
initial
begin
end

endmodule
