//-----------------------------------------------------------------------------
// File              : testcase2.sv
// Description       : Assembler code for test case 2 of the directed tests.
//                     This test exercises arithmetic and logical instructions.
// Pimrary Author    : Lewis Russell
// Other Contributers:
//------------------------------------------------------------------------------
32'h3C011234, // li     $1,      0x12340000
32'h34215678, // ori    $1,  $1, 0x5678
32'h3C020123, // li     $2,      0x01230000
32'h34424567, // ori    $2,  $2, 0x4567
32'h00221820, // add    $3,  $1, $2
32'h00222022, // sub    $4,  $1, $2
32'h20455500, // addi   $5,  $2, 0x5500
32'h00223024, // and    $6,  $1, $2
32'h30277654, // andi   $7,  $1, 0x7654
32'h00224025, // or     $8,  $1, $2
32'h00224826, // xor    $9,  $1, $2
32'h00225027, // nor   $10,  $1, $2
32'h382B5555, // xori  $11,  $1, 0x5555
32'h302CFFFF, // andi  $12,  $1, 0xFFFF
32'h718D6820, // clz   $13, $12
32'h000C7022, // sub   $14,  $0, $12
32'h71CF7821, // clo   $15, $14
32'h00228021, // addu  $16,  $1, $2
32'h00228823, // subu  $17,  $1, $2
32'h24525500, // addiu $18,  $2, 0x5500
32'h00000000, // nop
32'h00000000, // nop
32'h00000000, // nop
32'h00000000, // nop
32'h00000000  // nop
