//----------------------------------------
// File: PIPE_tb.sv
// Description: Pipeline registers testbench
// Primary Author: Jack Barnes
// Other Contributors:
// Notes: Full test coverage
//----------------------------------------
module PIPE_tb;

timeunit 10ns; timeprecision 100ps;
const int clk = 100;

PIPE PIPE0 (
);

//Initial conditions
initial
begin
end

//Testing procedure
initial
begin
end

endmodule
