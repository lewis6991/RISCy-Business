//------------------------------------------------------------------------------
// File              : mux.sv
// Description       : Standard 2:1 32-bit signal multiplexer
// Primary Author    : Dominic Murphy
// Other Contributors: Lewis Russell
// Notes             : - When sel is 0, Y = A. Else, Y = B.
//                     - Parameter n determines the bit width.
//------------------------------------------------------------------------------

module mux #(parameter n = 32)(
    input                Sel,
    input        [n-1:0] A  ,
                         B  ,
    output logic [n-1:0] Y
);

assign Y = Sel ? B : A;

endmodule
