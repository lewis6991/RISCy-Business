//-----------------------------------------------------------------------------
// File              : testcase4.sv
// Description       : Assembler code for test case 4 of the directed tests.
//                     This test exercises shift instructions.
// Pimrary Author    : Lewis Russell
// Other Contributers:
//------------------------------------------------------------------------------
32'h3C018005, // li    $1 ,      0x80050000
32'h34420004, // ori   $2 , $2 , 0x4
32'h00011943, // sra   $3 , $1 , 0x5
32'h00412007, // srav  $4 , $1 , $2
32'h00012940, // sll   $5 , $1 , 0x5
32'h00013142, // srl   $6 , $1 , 0x5
32'h00413804, // sllv  $7 , $1 , $2
32'h00414006, // srlv  $8 , $1 , $2
32'h0027480B, // movn  $9 , $1 , $7
32'h00C0500A, // movz  $10, $6 , $0
32'h0046582A, // slt   $11, $2 , $6
32'h284C0100, // slti  $12, $2 , 0x0100
32'h3C0D8800, // li    $13,      0x88000000
32'h002D702B, // sltu  $14, $1 , $13
32'h2D6F3200, // sltiu $15, $11, 0x3200
32'h00000000, // nop
32'h00000000, // nop
32'h00000000, // nop
32'h00000000, // nop
32'h00000000  // nop
