//------------------------------------------------------------------------------
// File              : branch_definition.sv
// Description       : Branch instruction codes
// Primary Author    : Dhanushan Raveendran
// Other Contributors: Lewis Russell, Ethan Bishop
// Notes             :
//------------------------------------------------------------------------------

`define BGEZ   6'b000001
`define BGEZAL 6'b010001
`define BLTZ   6'b000000
`define BLTZAL 6'b010000
