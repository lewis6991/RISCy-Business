//----------------------------------------
// File: FU_tb.sv
// Description: Data forwarding unit testbench
// Primary Author: Jack Barnes
// Other Contributors:
// Notes: Full test coverage
//----------------------------------------
module FU_tb;

timeunit 10ns; timeprecision 100ps;
const int clk = 100;

FU FU0 (
);

//Initial conditions
initial
begin
end

//Testing procedure
initial
begin
end

endmodule
