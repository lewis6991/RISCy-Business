//-----------------------------------------------------
// File: processor.sv
// Description: Top-level module for MIPS32 processor.
//-----------------------------------------------------

module processor(
    input logic Clock,
    input logic nReset
);

endmodule
