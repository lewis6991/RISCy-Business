//------------------------------------------------------------------------------
// File              : WB.sv
// Description       : Write Back pipeline stage
// Primary Author    : Dominic Murphy
// Other Contributors: Lewis Russell
// Notes             : - A very basic stage. Simple a mux, along with some
//                       control wires.
//                     - Warning: Names have no meaning yet, hence have been
//                       arbitrarily chosen.
//------------------------------------------------------------------------------

module WB(
    input        [31:0] Jack , 
                        Ethan,
    output logic [31:0] Lewis,
    output logic        Dhanu
);

    mux mux3(
        .Sel(UNKNOWN),
        .A  (Jack   ),
        .B  (Ethan  ),
        .Y  (Lewis  )
    );

endmodule
