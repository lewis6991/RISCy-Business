//----------------------------------------
// File: MEM_tb.sv
// Description: Memory testbench
// Primary Author: Jack Barnes
// Other Contributors:
// Notes: Full test coverage
//----------------------------------------
module MEM_tb;

timeunit 10ns; timeprecision 100ps;
const int clk = 100;

MEM MEM0 (
);

//Initial conditions
initial
begin
end

//Testing procedure
initial
begin
end

endmodule
