//----------------------------------------
// File: alu.sv
// Description: Arithmetic Logic Unit
// Primary Author: Ethan Bishop
// Other Contributors: Lewis Russell
//----------------------------------------

module alu(
    input        [31:0] A,
    input        [31:0] B,
    input        [4:0]  Shamt,
    input        [5:0]  ALUfunc,
    output logic [31:0] Out,
    output logic        En, C, Z, O, N
);

always_comb:
begin

    Out = 0;
    En = 1;
    C = 0;
    O = 0;
    N = Out[31];
    Z = (Out == 0);
    
    case (Func)
        ADD:
            begin
                {C, Out} = A + B;
                if (A[31] == B[31])
                    O = (A[31] ^ N);
            end
        ADDU:
            begin
                {C, Out} = A + B;
                O = C;
            end
        SUB:
            begin
                {C, Out} = A - B;
                if (A[31] == B[31])
                    O = (A[31] ^ N);
            end
        SUBU:
            begin
                {C, Out} = A - B;
                O = C;
            end
            
        SLL:
            Out = B << Shamt;
        SLLV:
            Out = B << A;
        SRA:
            Out = B >>> Shamt;
        SRAV:
            Out = B >>> A;
        SRL:
            Out = B >> Shamt;
        SRLV:
            Out = B >> A;

        AND:
            Out = A & B;
        NOR:
            Out = ~(A | B);
        OR:
            Out = A | B;
        XOR:
            Out = A ^ B;

        MOVN:
            begin
                Out = A;
                En = (B != 0);
            end
        MOVZ:
            begin
                Out = A;
                En = (B == 0);
            end
        
        SLT:
            if ((int)A < (int)B)
                Out = 1;
            else
                Out = 0;
        SLTU:
            if ((unsigned int)A < (unsigned int)B)
                Out = 1;
            else
                Out = 0;

        ALU_CLZ:
            case (A)
                32'b1???????????????????????????????: Out = 0;
                32'b01??????????????????????????????: Out = 1;
                32'b001?????????????????????????????: Out = 2;
                32'b0001????????????????????????????: Out = 3;
                32'b00001???????????????????????????: Out = 4;
                32'b000001??????????????????????????: Out = 5;
                32'b0000001?????????????????????????: Out = 6;
                32'b00000001????????????????????????: Out = 7;
                32'b000000001???????????????????????: Out = 8;
                32'b0000000001??????????????????????: Out = 9;
                32'b00000000001?????????????????????: Out = 10;
                32'b000000000001????????????????????: Out = 11;
                32'b0000000000001???????????????????: Out = 12;
                32'b00000000000001??????????????????: Out = 13;
                32'b000000000000001?????????????????: Out = 14;
                32'b0000000000000001????????????????: Out = 15;
                32'b00000000000000001???????????????: Out = 16;
                32'b000000000000000001??????????????: Out = 17;
                32'b0000000000000000001?????????????: Out = 18;
                32'b00000000000000000001????????????: Out = 19;
                32'b000000000000000000001???????????: Out = 20;
                32'b0000000000000000000001??????????: Out = 21;
                32'b00000000000000000000001?????????: Out = 22;
                32'b000000000000000000000001????????: Out = 23;
                32'b0000000000000000000000001???????: Out = 24;
                32'b00000000000000000000000001??????: Out = 25;
                32'b000000000000000000000000001?????: Out = 26;
                32'b0000000000000000000000000001????: Out = 27;
                32'b00000000000000000000000000001???: Out = 28;
                32'b000000000000000000000000000001??: Out = 29;
                32'b0000000000000000000000000000001?: Out = 30;
                32'b00000000000000000000000000000001: Out = 31;
                32'b00000000000000000000000000000000: Out = 32;
            endcase
            
        ALU_CLO:
            case (A)
                32'b0???????????????????????????????: Out = 0;
                32'b10??????????????????????????????: Out = 1;
                32'b110?????????????????????????????: Out = 2;
                32'b1110????????????????????????????: Out = 3;
                32'b11110???????????????????????????: Out = 4;
                32'b111110??????????????????????????: Out = 5;
                32'b1111110?????????????????????????: Out = 6;
                32'b11111110????????????????????????: Out = 7;
                32'b111111110???????????????????????: Out = 8;
                32'b1111111110??????????????????????: Out = 9;
                32'b11111111110?????????????????????: Out = 10;
                32'b111111111110????????????????????: Out = 11;
                32'b1111111111110???????????????????: Out = 12;
                32'b11111111111110??????????????????: Out = 13;
                32'b111111111111110?????????????????: Out = 14;
                32'b1111111111111110????????????????: Out = 15;
                32'b11111111111111110???????????????: Out = 16;
                32'b111111111111111110??????????????: Out = 17;
                32'b1111111111111111110?????????????: Out = 18;
                32'b11111111111111111110????????????: Out = 19;
                32'b111111111111111111110???????????: Out = 20;
                32'b1111111111111111111110??????????: Out = 21;
                32'b11111111111111111111110?????????: Out = 22;
                32'b111111111111111111111110????????: Out = 23;
                32'b1111111111111111111111110???????: Out = 24;
                32'b11111111111111111111111110??????: Out = 25;
                32'b111111111111111111111111110?????: Out = 26;
                32'b1111111111111111111111111110????: Out = 27;
                32'b11111111111111111111111111110???: Out = 28;
                32'b111111111111111111111111111110??: Out = 29;
                32'b1111111111111111111111111111110?: Out = 31;
                32'b11111111111111111111111111111110: Out = 31;
                32'b11111111111111111111111111111111: Out = 32;
            endcase
        
    endcase
    
end

endmodule
