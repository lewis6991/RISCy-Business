//---------------------------------------------
// File: Control.sv
// Description: Control module.
//---------------------------------------------

module control(
    input logic Clock,
    input logic nReset,
);

endmodule
