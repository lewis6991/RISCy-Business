//----------------------------------------
// File: EX_tb.sv
// Description: Execute testbench
// Primary Author: Jack Barnes
// Other Contributors:
// Notes: Full test coverage
//----------------------------------------
module EX_tb;

timeunit 10ns; timeprecision 100ps;
const int clk = 100;

EX EX0 (
);

//Initial conditions
initial
begin
end

//Testing procedure
initial
begin
end

endmodule
