//----------------------------------------
// File: control_tb.sv
// Description: Control testbench
// Primary Author: Jack Barnes
// Other Contributors:
// Notes: Full test coverage
//----------------------------------------
module control_tb;

timeunit 10ns; timeprecision 100ps;
const int clk = 100;

control control0 (
);

//Initial conditions
initial
begin
end

//Testing procedure
initial
begin
end

endmodule
