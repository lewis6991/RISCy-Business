//------------------------------------------------
// File: registers.sv
// Description: Register file module of 32x32-bit registers.
//------------------------------------------------

module registers(

);


endmodule
