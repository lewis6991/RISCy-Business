//----------------------------------------
// File: forwarding_unit_tb.sv
// Description: Data forwarding unit testbench
// Primary Author: Jack Barnes
// Other Contributors:
// Notes: Full test coverage
//----------------------------------------
module forwarding_unit_tb;

timeunit 10ns; timeprecision 100ps;
const int clk = 100;

forwarding_unit forwarding_unit0 (
);

//Initial conditions
initial
begin
end

//Testing procedure
initial
begin
end

endmodule
