//----------------------------------------
// File: alu.sv
// Description: Arithmetic Logic Unit
//----------------------------------------
module alu(
    input  logic [31:0] A   ,
    input  logic [31:0] B   ,
    output logic [31:0] Out ,
    input  logic [ 5:0] Func,
);


endmoudule
