//----------------------------------------
// File: WB_tb.sv
// Description: Write Back testbench
// Primary Author: Jack Barnes
// Other Contributors:
// Notes: Full test coverage
//----------------------------------------
module WB_tb;

timeunit 10ns; timeprecision 100ps;
const int clk = 100;

WB WB0 (
);

//Initial conditions
initial
begin
end

//Testing procedure
initial
begin
end

endmodule
