//------------------------------------------------------------------------------
// File              : BP.sv
// Description       : Branch prediction unit
// Primary Author    : -
// Other Contributors: 
// Notes             : Placeholder
//------------------------------------------------------------------------------

module BP(
    input        placeIn ,
    output logic placeOut
);

assign placeOut = placeIn;

endmodule
